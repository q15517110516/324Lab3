
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MUX IS
  PORT(    
  D0       : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
   D1        : IN STD_LOGIC_VECTOR(7 DOWNTO 0); 
   Y        : OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
   SEL     : IN  STD_LOGIC
      );
END ENTITY MUX;

ARCHITECTURE BEHAV OF MUX IS
BEGIN
    
         Y <= D0 when SEL='1' else  
              D1;    

 END ARCHITECTURE BEHAV;